module  FFT (
	input clk,
	input rst,
	input [15:0] fir_d, 
	input fir_valid, 
	output fftr_valid, 
	output ffti_valid, 
	output done,
	output [15:0] fft_d0
 	output [15:0] fft_d1, 
	output [15:0] fft_d2,
	output [15:0] fft_d3,
	output [15:0] fft_d4,
	output [15:0] fft_d5,
	output [15:0] fft_d6,
	output [15:0] fft_d7,
	output [15:0] fft_d8,
 	output [15:0] fft_d9,
	output [15:0] fft_d10,
	output [15:0] fft_d11,
	output [15:0] fft_d12,
	output [15:0] fft_d13,
	output [15:0] fft_d14,
	output [15:0] fft_d15
);

/////////////////////////////////
// Please write your code here //
/////////////////////////////////

endmodule