module BU(
	input signed [31:0] a,
	input signed [31:0] b,
	input signed [31:0] c,
	input signed [31:0] d,
	input signed [31:0] W_real,
	input signed [31:0] W_imag,
	
	output signed [31:0] result0_real,
	output signed [31:0] result0_imag,
	output signed [31:0] result1_real,
	output signed [31:0] result1_imag
);

/////////////////////////////////
// Please write your code here //
/////////////////////////////////

endmodule